
 
 
 

 



window new WaveWindow  -name  "Waves for BMG Example Design"
waveform  using  "Waves for BMG Example Design"


      waveform add -signals /startpage_tb/status
      waveform add -signals /startpage_tb/startpage_synth_inst/bmg_port/CLKA
      waveform add -signals /startpage_tb/startpage_synth_inst/bmg_port/ADDRA
      waveform add -signals /startpage_tb/startpage_synth_inst/bmg_port/DINA
      waveform add -signals /startpage_tb/startpage_synth_inst/bmg_port/WEA
      waveform add -signals /startpage_tb/startpage_synth_inst/bmg_port/DOUTA
console submit -using simulator -wait no "run"
