`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:38:25 12/31/2019 
// Design Name: 
// Module Name:    show_back 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module show_back(
			input ad;
			input clk;
			output col;
    );
		always@(posedge clk)begin
			case(ad)
				
		
		
		end

endmodule
